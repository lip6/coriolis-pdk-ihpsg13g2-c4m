.subckt tie_diff vdd vss
.ends tie_diff
