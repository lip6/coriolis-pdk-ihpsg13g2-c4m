.subckt or21nand_x0 vdd vss nq i0 i1 i2
Xi0_nmos _net0 i0 vss vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi0_pmos vdd i0 _net1 vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi1_nmos vss i1 _net0 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi1_pmos _net1 i1 nq vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi2_nmos _net0 i2 nq vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi2_pmos nq i2 vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
.ends or21nand_x0
