.subckt dff_x1 vdd vss i clk q
Xclk_nmos _clk_n clk vss vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xclk_pmos _clk_n clk vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xclk_n_nmos0 vss _clk_n _clk_buf vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xclk_n_pmos0 vdd _clk_n _clk_buf vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi_nmos _u i vss vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi_pmos _u i vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xu_nmos vss _u _net0 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xu_pmos vdd _u _net1 vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xclk_n_nmos1 _net0 _clk_n _dff_m vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xclk_buf_pmos0 _net1 _clk_buf _dff_m vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xclk_buf_nmos0 _dff_m _clk_buf _net2 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xclk_n_pmos1 _dff_m _clk_n _net3 vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xy_nmos _net2 _y vss vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xy_pmos _net3 _y vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xdff_m_nmos vss _dff_m _y vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xdff_m_pmos vdd _dff_m _y vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xclk_buf_nmos1 _y _clk_buf _dff_s vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xclk_n_pmos2 _y _clk_n _dff_s vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xclk_n_nmos2 _dff_s _clk_n _net4 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xclk_buf_pmos1 _dff_s _clk_buf _net5 vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xq_nmos _net4 q vss vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xq_pmos _net5 q vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xdff_s_nmos vss _dff_s q vss sg13_lv_nmos l=1.3e-07 w=9.4e-07
Xdff_s_pmos vdd _dff_s q vdd sg13_lv_pmos l=1.3e-07 w=9.8e-07
.ends dff_x1
