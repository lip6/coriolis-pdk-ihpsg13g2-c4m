.subckt nor3_x1 vdd vss nq i0 i1 i2
Xi0_nmos vss i0 nq vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi0_pmos vdd i0 _net0 vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi1_nmos nq i1 vss vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi1_pmos _net0 i1 _net1 vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi2_nmos vss i2 nq vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi2_pmos _net1 i2 nq vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
.ends nor3_x1
