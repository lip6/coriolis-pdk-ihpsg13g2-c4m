.subckt tie_poly_w4 vdd vss
.ends tie_poly_w4
