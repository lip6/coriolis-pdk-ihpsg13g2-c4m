.subckt tie_diff_w2 vdd vss
.ends tie_diff_w2
