.subckt or2_x1 vdd vss q i0 i1
Xi0_nmos vss i0 nq vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi0_pmos nq i0 _net0 vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi1_nmos nq i1 vss vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi1_pmos _net0 i1 vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xn_pd vss nq q vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xq_pu vdd nq q vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
.ends or2_x1
