.subckt nand2_x1 vdd vss nq i0 i1
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi1_nmos _net0 i1 nq vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
.ends nand2_x1
