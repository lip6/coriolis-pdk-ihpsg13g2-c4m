.subckt diode_w1 vdd vss i
.ends diode_w1
