.subckt tie_poly_w2 vdd vss
.ends tie_poly_w2
