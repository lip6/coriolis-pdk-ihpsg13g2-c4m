.subckt fill_w4 vdd vss
.ends fill_w4
