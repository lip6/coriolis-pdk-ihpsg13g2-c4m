.subckt nand3_x1 vdd vss nq i0 i1 i2
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi1_nmos _net0 i1 _net1 vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi2_nmos _net1 i2 nq vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi2_pmos vdd i2 nq vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
.ends nand3_x1
