.subckt fill_w2 vdd vss
.ends fill_w2
