.subckt nand4_x0 vdd vss nq i0 i1 i2 i3
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi1_nmos _net0 i1 _net1 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi2_nmos _net1 i2 _net2 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi2_pmos vdd i2 nq vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi3_nmos _net2 i3 nq vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi3_pmos nq i3 vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
.ends nand4_x0
