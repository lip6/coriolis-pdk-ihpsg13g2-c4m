.subckt and21nor_x1 vdd vss nq i0 i1 i2
Xi0_nmos vss i0 _net1 vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi0_pmos _net0 i0 vdd vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi1_nmos _net1 i1 nq vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi1_pmos vdd i1 _net0 vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
Xi2_nmos nq i2 vss vss sg13_lv_nmos l=1.3e-07 w=1.66e-06
Xi2_pmos _net0 i2 nq vdd sg13_lv_pmos l=1.3e-07 w=1.7e-06
.ends and21nor_x1
