.subckt tie_diff_w4 vdd vss
.ends tie_diff_w4
