.subckt nsnrlatch_x1 vdd vss nset nrst q nq
Xnset_nmos q nset _net0 vss sg13_lv_nmos l=1.3e-07 w=1.48e-06
Xnset_pmos vdd nset q vdd sg13_lv_pmos l=1.3e-07 w=1.52e-06
Xnq_nmos _net0 nq vss vss sg13_lv_nmos l=1.3e-07 w=1.48e-06
Xnq_pmos q nq vdd vdd sg13_lv_pmos l=1.3e-07 w=1.52e-06
Xq_nmos vss q _net1 vss sg13_lv_nmos l=1.3e-07 w=1.48e-06
Xq_pmos vdd q nq vdd sg13_lv_pmos l=1.3e-07 w=1.52e-06
Xnrst_nmos _net1 nrst nq vss sg13_lv_nmos l=1.3e-07 w=1.48e-06
Xnrst_pmos nq nrst vdd vdd sg13_lv_pmos l=1.3e-07 w=1.52e-06
.ends nsnrlatch_x1
