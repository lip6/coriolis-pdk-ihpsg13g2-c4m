.subckt nand3_x0 vdd vss nq i0 i1 i2
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi1_nmos _net0 i1 _net1 vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
Xi2_nmos _net1 i2 nq vss sg13_lv_nmos l=1.3e-07 w=7.8e-07
Xi2_pmos vdd i2 nq vdd sg13_lv_pmos l=1.3e-07 w=7.8e-07
.ends nand3_x0
